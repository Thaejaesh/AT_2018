library verilog;
use verilog.vl_types.all;
entity MATRIX_MULTIPLIER_v_unit is
end MATRIX_MULTIPLIER_v_unit;
