library verilog;
use verilog.vl_types.all;
entity Milestone_2_v_unit is
end Milestone_2_v_unit;
