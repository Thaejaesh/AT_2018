library verilog;
use verilog.vl_types.all;
entity WS_v_unit is
end WS_v_unit;
