library verilog;
use verilog.vl_types.all;
entity MATRIX_MULT_v_unit is
end MATRIX_MULT_v_unit;
