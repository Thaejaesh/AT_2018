library verilog;
use verilog.vl_types.all;
entity FS_v_unit is
end FS_v_unit;
