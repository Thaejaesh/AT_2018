library verilog;
use verilog.vl_types.all;
entity Milestone_3_v_unit is
end Milestone_3_v_unit;
